module counter(
